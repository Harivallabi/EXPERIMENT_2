module mux(d,s,y);
input[7:0]d;
input[2:0]s;
output y;
wire w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11;
not g1 (w1,s[2]);
not g2(w2,s[1]);
not g3(w3,s[0]);
and g4(w4,w1,w2,w3,d[0]);
and g5(w5,w1,w2,s[0],d[1]);
and g6(w6,w1,w3,s[1],d[2]);
and g7(w7,w1,s[1],s[0],d[3]);
and g8(w8,w2,w3,s[2],d[4]);
and g9(w9,w2,s[2],s[0],d[5]);
and g10(w10,w3,s[1],s[2],d[6]);
and g11(w11,s[0],s[1],s[2],d[7]);
or g12(y,w4,w5,w6,w7,w8,w9,w10,w11);
endmodule
